`timescale 1ns / 1ps
module Word(
	output reg	[679:0]	word	,			//��ģ������
	input			[5:0]		choose			//��ģ����	
    );
	 
always @(*) begin
	Word_Choose(choose);						//������ģ��ѡ������
	end

task Word_Choose;
	input	[5:0] d;
	begin
		case (d)
			0: word = 680'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;			1: word = 680'h00080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000060000000000040000000000000;			2: word = 680'h001C1800000000600000003000000000070180000000400C00000001000000000000000000000000000000000000000000000000000000000000000000180000000020000000000030000000000060000000600000;			3: word = 680'h001C0C000000003000000038000030000300E0000040600F00000000C000000000000000000000000000000000000000000000000000000000000000001E000030003800006000001C000000040070000000380000;			4: word = 680'h00180E000000003800000031FFFFF8000300C0200060300E000C0C00E0000000000000000000000000000000000000000000000000000000000000000038000030001C0001F000001C0000000E00E00000001C0000;			5: word = 680'h003806000000001C00000030C06000000300C0700030381C000FFE006000000000000000000003000000000000000000000000000000000000000000003F000030001C218FE000000E00001FFE00D00000001C0000;			6: word = 680'h00300400C000001C000000300060003FFFFFFFF800383818000C1C406020000007F0FC003000FF000030000000000000000001F8801F807FF8000F880071C00030000871F00000000C0000000C01D0000200080020;			7: word = 680'h007FFFFFE000001800000C300060001C0300C000001C1C18000C18404070000001C030007800070000780000000000000000060F8030C01C0E0038780070E000301FFFF9C00002000C0020000C0188000200000060;			8: word = 680'h00E00C000002000000600F30006000000300C000001C1830000C18FFFFF0000001C0200078000700007800000000000000000C0380E0701C030060180060780030080080C0000200000070020C038C0003FFFFFFF0;			9: word = 680'h00E00C000003FFFFFFF00E30006000000300C000001C1820000C10C00040000000E0600030000700003000000000000000001C0180C0301C0380C01800C03C20300101C0C00003FFFFFFF8078C03040006000000E0;			10:word = 680'h01E00C000002000000780E30006000000300C00002080040100C31C00080000000E04000000007000000000000000000000038018180181C01C1C00C00C01C38300181C0C0000600000070060C0606000600000080;			11:word = 680'h03600C030006000000C00E30806020000300800002000040300C21C00080000000704000000007000000000000000000000038008380181C01C1800401800C303000C180C00006080600C0060C0603000E00000500;			12:word = 680'h067FFFFF8006000001800630FFFFF8018000000007FFFFFFF80C200000000000007080000000070000000000000000000000380083801C1C01C38004030000303000E300C0000E06078080060C0C03800E00000E00;			13:word = 680'h0C600C00000E000001000630C0603000E000020006000000700C400006000000003080000000070000000000000000000000380003000C1C01C38000030000303000E200C0000E07870100061C1801C001FFFFFF00;			14:word = 680'h08600C00000C000002000630C06030007030078006000000600C403FFF0000000039800030000700003000400000000000003C0003000C1C01C300000700403030004218C0300C0387000006181000F00000700000;			15:word = 680'h10600C020000000000C00630C0603000313FFF800E000000800C4000000000000039000FF00007000FF007C7C03F9F8000001E0007000E1C01C7000005FFE0303000043CC0780001C70000061820037C0000E00000;			16:word = 680'h207FFFFF0000000001E00630C0603000323003000E000019000C200000000000001F000070000700007001C8E00F060000001F0007000E1C0387000009807030301FFFFEFFFC000187000006185FFFB00001802000;			17:word = 680'h00600C00000FFFFFFFF00630C0603010023003001CFFFFF8000C100000000000001E000070000700007001D06007040000000FC007000E1C030700001980603030000C00C18000808700000E188E00000003001800;			18:word = 680'h00600C000000001800000630C060300C023003000040003C000C180000400000000E000070000700007001E070070C00000003F007000E1C0E0700002180E03030000C00C18000600700000C190000000006001C00;			19:word = 680'h00600C008000001800000630C06030060430030000000070000C0C0000E00000000E000070000700007001C070039800000000FC07000E1FFC0700000180E03030000C00C18000780600000C1B0000000018000E00;			20:word = 680'h00600C01C000001800000630C060300704300700000000C0000C0CFFFFF07FFFC00F000070000700007001C0700390000000003F07000E1C000700000180E03030000C00C180003C0600000FFF8100C000F0000700;			21:word = 680'h007FFFFFE000001800000630C06030038830070000000300000C060630000000000F000070000700007001C07001F0000000000F87000E1C000700000180E03030000C31C180001C06000004032180E0007FFFFF00;			22:word = 680'h006010000000001800000630C06030030830070000001600000C060630000000000B800070000700007001C07001E0000000000787000E1C000700000180C030300FFFF9C180001C06000000031080E0007E000300;			23:word = 680'h00601C000000001800000E30C06030001830060000001C00200C0606300000000013800070000700007001C07000E00000000003C7000E1C000700000180C03030000C01818000080E0030000310C0C00000180300;			24:word = 680'h000018001000001800000E30C06030001030060000001C00700C0606300000000013C00070000700007001C07000F00000000001C3000C1C000700000180C03030000C01818000000E0078000318E1C000001C0000;			25:word = 680'h000018003800001800000E60C0603000303086003FFFFFFFF80D0E06300000000021C00070000700007001C07000F00000002001C3800C1C00038004018FC03030010D0181801FFFFFFFFC000F1861800000180000;			26:word = 680'h3FFFFFFFFC00001800000860C060300020307E0018001C00000CFC0E300000000021E00070000700007001C07001380000002001C3801C1C00038004018784203003CC81818000000C000001F60C71800000180600;			27:word = 680'h0000F9000000001800000060C060300060301C2000001C00000C380C301000000060E00070000700007001C07003380000003001C1801C1C000380080183040030038CE1818000001C00003F060C71000000180F00;			28:word = 680'h0001D98000000018000000C0C063F007E030081000001C00000C200C301000000040E00070000700007001C070021C0000001001C180181C000180080180040030030C73018000001C000038060C730000FFFFFF80;			29:word = 680'h000398C000000018000000C0C060E001C030001000001C00000C001C3010000000C0700070000700007001C070041E000000180380C0301C0001C0100180040030060C33018000003B800010060C62000000180000;			30:word = 680'h0006186000000018000001808060C000C030003000001C00000C0018301000000080700070000700007001C0700C0E0000001C030060701C0000E0300180040030060C320180000070F00000060C02000000180000;			31:word = 680'h001C1838000000180000018000600000C030003000001C00000C0038301000000180780070000700007001C0701C0F0000001E0E0030C01C0000704001800400300C0C2601800000E03E0000060C06000000180000;			32:word = 680'h0038181C000000180000030000600000C030003800001C00000C00703010000007E0FE0FFF80FFF80FFF87F1FC7E3FC0000011FC001F807F00001F800180060030080C0C01800001C01F80000E0004000000180000;			33:word = 680'h00E0180F80000E380000020000600000C038007800001C00000C00E0383800000000000000000000000000000000000000000000000000000000000001800F0070101C08018000038007C0039C0004100000180030;			34:word = 680'h01801803FC0003F80000040000600000C01FFFF00003FC00000C01801FF800000000000000000000000000000000000000000000000000000000000001FFFE0FF020FC100180000E0003C000FC0008380000180078;			35:word = 680'h06001800F80000F00000080000600000C00000000000F800000C03001FF0000000000000000000000000000000000000000000000000000000000000007FF803E0003820018000780001C00078FFFFFC1FFFFFFFFC;			36:word = 680'h18001800300000700000100000600000C000000000007000000C1C00000000000000000000000000000000000000000000000000000000000000000000000000C0003040038003C00000C000200000000000000000;			37:word = 680'h200010000000004000002000004000000000000000002000000800000000000000000000000000000000000000000000000000000000000000000000000000000000008002001C0000000000000000000000000000;			38:word = 680'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;			39:word = 680'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			endcase
		end
	endtask

endmodule
